/* Hello World in Verilog. */

module main;

 initial
   begin
     $display("Hello, World");
     $finish ;
   end

 endmodule
